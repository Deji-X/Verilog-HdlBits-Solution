module top_module(
  input  [99:0]  in,
  output [99:0] out,
);
/* integer w;
    always @ (in) begin 
        for (w=0; w<100; w=w+1) begin
            out[99-w] = in[w];
        end        
    end
*/  

endmodule
