// Tb/tb1

module top_module(
  output reg A,
  output reg B
);

  initial begin

  end

endmodule
