//Tb/tff

module top_module(
  
);

endmodule
