module top_module(
  input clk,
  input [31:0] in,
  output [31:0] out
);

  

endmodule
