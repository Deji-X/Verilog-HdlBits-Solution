// Adder100

module top_module(
  input [99:0] a, b,
  input cin,
  output cout,
  output [99:0] sum
);

  wire 
  //This a 100 bit number, I am not going to write a function for 100 bits each,
  //hence, genvar i...generate.

  

endmodule
