// Adder100

module top_module(
  
);

endmodule
