// sim/circuit

module top_module(
  input clock,
  input a,
  output p,
  output q
);

  

endmodule
