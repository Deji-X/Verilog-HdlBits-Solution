module top_module(
  input clk,
  input [7:0] in,
  input [7:0] pedge
);

endmodule
