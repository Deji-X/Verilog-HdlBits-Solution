module top_module( input in, output out);
  assign out = ~in;
  // ~ is the bitwise function for "NOT"
  // | is the bitwise function for "OR"
  // & is the bitwise function for "AND"
endmodule
