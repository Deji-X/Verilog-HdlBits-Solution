// Tb/tb2
module top_module(
  
);

endmodule
