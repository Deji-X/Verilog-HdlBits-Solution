module top_mod(
  input clk,
  input d,
  output q
);
  wire clk
