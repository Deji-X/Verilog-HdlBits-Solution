module top_module(
  input clk,
  input areset, //Asynchronous reset to state B
  input in,
  output out
);

  parameter A=0, B=1;
  reg state, next_state;

  always @(*) begin  //This is a combinational always block
      //  State transition logic
  end

  always @ (posedge clk, posedge reset) begin  // This is a sequential always block
    // State flip-flops with asynchronous reset
  end

  // Output logic
  // assign out = (state == ....);

endmodule
