module top_module(
  input clk,
  input w, R, E, L,
  output Q
);

  wire 
